library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cpu is
end cpu;

architecture cpu of cpu is
begin
end cpu;
